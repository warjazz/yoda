module control(
input clk_100,
input BTNL,
input BTNR,
input BTNN,
input BTNS,
input BTNC)

parameter N = 'd12;
reg []

